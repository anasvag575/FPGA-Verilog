`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: ---
// Engineer: Vagenas Anastasis 2496
//
// Create Date:    20:10:01 10/12/2019
// Design Name:  -----
// Module Name:   VRAM
// Project Name: VGA Driver Lab03 Project
// Target Devices: FPGA Spartan 3E
// Tool versions: -----
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////
module vram_unit (clk,addr,r_pixel,g_pixel,b_pixel);

input clk;
input [13:0] addr;
output r_pixel,g_pixel,b_pixel;

RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_02(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_03(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_05(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_06(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_08(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_09(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0C(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_0E(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_0F(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_11(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_12(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_14(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_15(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_17(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_18(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_1A(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_1B(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_1D(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_1E(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      // Address 8192 to 12287
      .INIT_20(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_21(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_23(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_24(256'hFFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00FFFF00FFFF00FFFF),
      .INIT_25(256'h0000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00),
      .INIT_26(256'h00F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F0),
      .INIT_27(256'hFFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F000),
      .INIT_28(256'h0000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00),
      .INIT_29(256'h00F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F0),
      .INIT_2A(256'hFFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F000),
      .INIT_2B(256'h0000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00),
      .INIT_2C(256'h00F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F0),
      .INIT_2D(256'hFFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F000),
      .INIT_2E(256'h0000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F00000FFFF00FFFF00),
      .INIT_2F(256'h00F00000F00000F00000FFFF00FFFF00FFFF00FFFF00F00000F00000F00000F0),
   ) red_vram (
      .DO(r_pixel),       // 1-bit Data Output
      .ADDR(addr),       // 14-bit Address Input
      .CLK(clk),        // Clock
      .EN(1'b1),        // RAM Enable Input
		.SSR(1'b0) ,      // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

	RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_02(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_03(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_05(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_06(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_08(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_09(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_0B(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_0C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_11(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_12(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_14(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_15(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_17(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_18(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_1A(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_1B(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_1D(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_1E(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      // Address 8192 to 12287
      .INIT_20(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_21(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_23(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_24(256'h0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF),
      .INIT_25(256'h000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F),
      .INIT_26(256'h0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00),
      .INIT_27(256'h0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF),
      .INIT_28(256'h000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F),
      .INIT_29(256'h0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00),
      .INIT_2A(256'h0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF),
      .INIT_2B(256'h000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F),
      .INIT_2C(256'h0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00),
      .INIT_2D(256'h0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF),
      .INIT_2E(256'h000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00000F00000F0FFF0F),
      .INIT_2F(256'h0F00000F00000F00000F00000F0FFF0F0FFF0F0FFF0F0FFF0F00000F00000F00)
   ) green_vram (
      .DO(g_pixel),       // 1-bit Data Output
      .ADDR(addr),       // 14-bit Address Input
      .CLK(clk),        // Clock
      .EN(1'b1),        // RAM Enable Input
		.SSR(1'b0) ,      // Synchronous Set/Reset Input
      .WE(1'b0)       // Write Enable Input
   );

	RAMB16_S1 #(
      .INIT(1'b0),  // Value of output RAM registers at startup
      .SRVAL(1'b0), // Output value upon SSR assertion
      .WRITE_MODE("READ_FIRST"), // WRITE_FIRST, READ_FIRST or NO_CHANGE

      // The forllowing INIT_xx declarations specify the initial contents of the RAM
      // Address 0 to 4095
      .INIT_00(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_01(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_02(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_03(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_04(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_05(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_06(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_07(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_08(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_09(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0A(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_0B(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_0C(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_0D(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_0E(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_0F(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 4096 to 8191
      .INIT_10(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_11(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_12(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_13(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_14(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_15(256'hFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_16(256'h00000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFF),
      .INIT_17(256'h000000000000000000000000FFFFFFFFFFFFFFFFFFFFFFFF0000000000000000),
      .INIT_18(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_19(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1A(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1B(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1C(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1D(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1E(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_1F(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      // Address 8192 to 12287
      .INIT_20(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_21(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_22(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_23(256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF),
      .INIT_24(256'h0FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFF),
      .INIT_25(256'h00F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF0),
      .INIT_26(256'hF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F000),
      .INIT_27(256'h0FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFF),
      .INIT_28(256'h00F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF0),
      .INIT_29(256'hF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F000),
      .INIT_2A(256'h0FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFF),
      .INIT_2B(256'h00F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF0),
      .INIT_2C(256'hF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F000),
      .INIT_2D(256'h0FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFF),
      .INIT_2E(256'h00F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F00000F00000F00FFFF0),
      .INIT_2F(256'hF00000F00000F00000F00000F00FFFF00FFFF00FFFF00FFFF00000F00000F000)
   ) blue_vram (
      .DO(b_pixel),       // 1-bit Data Output
      .ADDR(addr),       // 14-bit Address Input
      .CLK(clk),        // Clock
      .EN(1'b1),       // RAM Enable Input
      .WE(1'b0)       // Write Enable Input
   );

endmodule
